library verilog;
use verilog.vl_types.all;
entity counter_vlg_tst is
end counter_vlg_tst;
